/************************************************/
/* Image Processor                              */
/*                                              */
/************************************************/

