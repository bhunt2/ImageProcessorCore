/************************************************/
/* Image Processor                              */
/*                                              */
/************************************************/

import ImageProcessingPkg::*;

module ImageProcessor(
	input clk,
	input rst,
	input pixel_t pixelA,
	input pixel_t pixelB,
	input opcodes_t opcode,
	output  result
);

	// Registers for pulling in and buffering data
	reg [

    // Bring in the 
    always_comb begin
		
    end

endmodule
