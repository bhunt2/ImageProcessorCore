import CellProcessingPkg::cellDepth;
import CellProcessingPkg::opCodeWidth;

// Interface
interface cellProcessor_int(input logic clk, rst);
    logic [cellDepth - 1:0] 		cellA;
    logic [cellDepth - 1:0] 		cellB;
    CellProcessingPkg::userInput_t  userInputA;
    logic [opCodeWidth - 1:0]		opcode;
    CellProcessingPkg::pixel_t		processedPixel;
    
    modport cellPorts ( input  clk,
                        input  rst,
                        input  cellA,
                        input  cellB,
                        input  userInputA,
                        input  opcode,
                        output processedPixel
                      );
                      
    modport imagePorts ( output cellA,
                         output cellB,
                         output userInputA,
                         output opcode
                       );
                       
endinterface